module fonts

// fonts - simple fonts for drawing on a canvas

// A very simple bitmap font...
// Stolen from https://github.com/mikaelpatel/Arduino-LCD/blob/master/src/Driver/PCD8544.h#L304 with minor tweaks
// Only does ASCII chars 32..127 in a 5x7 font in a 6x8 cell

pub const (
	simple_font             = [
		0x00,
		0x00,
		0x00,
		0x00,
		0x00,
		0x00,
		0x00,
		0x5F,
		0x00,
		0x00,
		0x00,
		0x07,
		0x00,
		0x07,
		0x00,
		0x14,
		0x7F,
		0x14,
		0x7F,
		0x14,
		0x24,
		0x2A,
		0x7F,
		0x2A,
		0x12,
		0x23,
		0x13,
		0x08,
		0x64,
		0x62,
		0x36,
		0x49,
		0x56,
		0x20,
		0x50,
		0x00,
		0x08,
		0x07,
		0x03,
		0x00,
		0x00,
		0x1C,
		0x22,
		0x41,
		0x00,
		0x00,
		0x41,
		0x22,
		0x1C,
		0x00,
		0x2A,
		0x1C,
		0x7F,
		0x1C,
		0x2A,
		0x08,
		0x08,
		0x3E,
		0x08,
		0x08,
		0x00,
		0x80,
		0x70,
		0x30,
		0x00,
		0x08,
		0x08,
		0x08,
		0x08,
		0x08,
		0x00,
		0x00,
		0x60,
		0x60,
		0x00,
		0x20,
		0x10,
		0x08,
		0x04,
		0x02,
		0x3E,
		0x51,
		0x49,
		0x45,
		0x3E,
		0x00,
		0x42,
		0x7F,
		0x40,
		0x00,
		0x72,
		0x49,
		0x49,
		0x49,
		0x46,
		0x21,
		0x41,
		0x49,
		0x4D,
		0x33,
		0x18,
		0x14,
		0x12,
		0x7F,
		0x10,
		0x27,
		0x45,
		0x45,
		0x45,
		0x39,
		0x3C,
		0x4A,
		0x49,
		0x49,
		0x31,
		0x41,
		0x21,
		0x11,
		0x09,
		0x07,
		0x36,
		0x49,
		0x49,
		0x49,
		0x36,
		0x46,
		0x49,
		0x49,
		0x29,
		0x1E,
		0x00,
		0x00,
		0x14,
		0x00,
		0x00,
		0x00,
		0x40,
		0x34,
		0x00,
		0x00,
		0x00,
		0x08,
		0x14,
		0x22,
		0x41,
		0x14,
		0x14,
		0x14,
		0x14,
		0x14,
		0x00,
		0x41,
		0x22,
		0x14,
		0x08,
		0x02,
		0x01,
		0x59,
		0x09,
		0x06,
		0x3E,
		0x41,
		0x5D,
		0x59,
		0x4E,
		0x7C,
		0x12,
		0x11,
		0x12,
		0x7C,
		0x7F,
		0x49,
		0x49,
		0x49,
		0x36,
		0x3E,
		0x41,
		0x41,
		0x41,
		0x22,
		0x7F,
		0x41,
		0x41,
		0x41,
		0x3E,
		0x7F,
		0x49,
		0x49,
		0x49,
		0x41,
		0x7F,
		0x09,
		0x09,
		0x09,
		0x01,
		0x3E,
		0x41,
		0x41,
		0x51,
		0x73,
		0x7F,
		0x08,
		0x08,
		0x08,
		0x7F,
		0x00,
		0x41,
		0x7F,
		0x41,
		0x00,
		0x20,
		0x40,
		0x41,
		0x3F,
		0x01,
		0x7F,
		0x08,
		0x14,
		0x22,
		0x41,
		0x7F,
		0x40,
		0x40,
		0x40,
		0x40,
		0x7F,
		0x02,
		0x1C,
		0x02,
		0x7F,
		0x7F,
		0x04,
		0x08,
		0x10,
		0x7F,
		0x3E,
		0x41,
		0x41,
		0x41,
		0x3E,
		0x7F,
		0x09,
		0x09,
		0x09,
		0x06,
		0x3E,
		0x41,
		0x51,
		0x21,
		0x5E,
		0x7F,
		0x09,
		0x19,
		0x29,
		0x46,
		0x26,
		0x49,
		0x49,
		0x49,
		0x32,
		0x03,
		0x01,
		0x7F,
		0x01,
		0x03,
		0x3F,
		0x40,
		0x40,
		0x40,
		0x3F,
		0x1F,
		0x20,
		0x40,
		0x20,
		0x1F,
		0x3F,
		0x40,
		0x38,
		0x40,
		0x3F,
		0x63,
		0x14,
		0x08,
		0x14,
		0x63,
		0x03,
		0x04,
		0x78,
		0x04,
		0x03,
		0x61,
		0x59,
		0x49,
		0x4D,
		0x43,
		0x00,
		0x7F,
		0x41,
		0x41,
		0x41,
		0x02,
		0x04,
		0x08,
		0x10,
		0x20,
		0x00,
		0x41,
		0x41,
		0x41,
		0x7F,
		0x04,
		0x02,
		0x01,
		0x02,
		0x04,
		0x40,
		0x40,
		0x40,
		0x40,
		0x40,
		0x00,
		0x03,
		0x07,
		0x08,
		0x00,
		0x20,
		0x54,
		0x54,
		0x78,
		0x40,
		0x7F,
		0x28,
		0x44,
		0x44,
		0x38,
		0x38,
		0x44,
		0x44,
		0x44,
		0x28,
		0x38,
		0x44,
		0x44,
		0x28,
		0x7F,
		0x38,
		0x54,
		0x54,
		0x54,
		0x18,
		0x00,
		0x08,
		0x7E,
		0x09,
		0x02,
		0x18,
		0xA4,
		0xA4,
		0x9C,
		0x78,
		0x7F,
		0x08,
		0x04,
		0x04,
		0x78,
		0x00,
		0x44,
		0x7D,
		0x40,
		0x00,
		0x20,
		0x40,
		0x40,
		0x3D,
		0x00,
		0x7F,
		0x10,
		0x28,
		0x44,
		0x00,
		0x00,
		0x41,
		0x7F,
		0x40,
		0x00,
		0x7C,
		0x04,
		0x78,
		0x04,
		0x78,
		0x7C,
		0x08,
		0x04,
		0x04,
		0x78,
		0x38,
		0x44,
		0x44,
		0x44,
		0x38,
		0xFC,
		0x18,
		0x24,
		0x24,
		0x18,
		0x18,
		0x24,
		0x24,
		0x18,
		0xFC,
		0x7C,
		0x08,
		0x04,
		0x04,
		0x08,
		0x48,
		0x54,
		0x54,
		0x54,
		0x24,
		0x04,
		0x04,
		0x3F,
		0x44,
		0x24,
		0x3C,
		0x40,
		0x40,
		0x20,
		0x7C,
		0x1C,
		0x20,
		0x40,
		0x20,
		0x1C,
		0x3C,
		0x40,
		0x30,
		0x40,
		0x3C,
		0x44,
		0x28,
		0x10,
		0x28,
		0x44,
		0x0C,
		0x90,
		0x90,
		0x90,
		0x7C,
		0x44,
		0x64,
		0x54,
		0x4C,
		0x44,
		0x00,
		0x08,
		0x36,
		0x41,
		0x00,
		0x00,
		0x00,
		0x7F,
		0x00,
		0x00,
		0x00,
		0x41,
		0x36,
		0x08,
		0x00,
		0x02,
		0x01,
		0x02,
		0x04,
		0x02,
		0x3C,
		0x26,
		0x23,
		0x26,
		0x3C,
	]
	simple_font_char_height = 7
	simple_font_char_width  = 5
)
